`define DATA_WIDTH     16
`define INST_WIDTH     64

`define PORTAWIDTH     30
`define PORTBWIDTH     18
`define PORTCWIDTH     48
`define PORTPWIDTH     48

`define REG_ADDR_WIDTH  8
`define DM_ADDR_WIDTH 	8
`define IM_ADDR_WIDTH 	8