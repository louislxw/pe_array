`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10.06.2020 17:00:46
// Design Name: 
// Module Name: tb_data_mem
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
`include "parameters.vh"

module tb_data_mem;

    // Inputs
    reg clk; 
    reg rst;
    reg wea; 
    reg web;
    reg [`DATA_WIDTH*2-1:0] dina;
    reg [`DATA_WIDTH*2-1:0] dinb;
    reg wben;
    reg rden;
    reg inst_v;
    reg [`INST_WIDTH-1:0] inst;
    
    // Outputs
    wire [`DATA_WIDTH*2-1:0] douta;
    wire [`DATA_WIDTH*2-1:0] doutb;


    // Instantiate the Unit Under Test (UUT)
    data_mem DMEM(
    .clk(clk), 
    .rst(rst), 
    .wea(wea), 
    .web(web),
    .dina(dina), 
    .dinb(dinb),
    .wben(wben),
    .rden(rden), 
    .inst_v(inst_v),
    .inst(inst), 
    .douta(douta),
    .doutb(doutb)
    );

    parameter PERIOD = 20;

    always begin
        clk = 1'b0;
        #(PERIOD/2) clk = 1'b1;
        #(PERIOD/2);
    end
    
    integer cycle;
    
    initial cycle = 0;
    always @(posedge clk)
        cycle = cycle + 1;
    
    initial begin
        // Initialize Inputs
        clk = 0;
        rst = 0;
        wea = 0;
        web = 0;
        dina = 0; 
        dinb = 0;
        wben = 0;
        rden = 0;
        inst_v = 0;
        inst = 0;
        
        // Wait 100 ns for global reset to finish
        rst = 1;
        #100;
        
        // Add stimulus here
        #20; wea = 0; rst = 0; 
		#20; wea = 0;  
		#20; wea = 0; 
		#20; wea = 0; 
        // wea or rden is aligned with inst; 1 cycle ahead of wdata 
        #20; wea = 0;                 
		#20; wea = 1; dina = 32'h0004_0002; // 4 + j*2 
		#20; wea = 1; dina = 32'h0003_0001; // 3 + j*1 
		#20; wea = 1; dina = 32'h0008_0006; // 8 + j*6 
		#20; wea = 1; dina = 32'h0007_0005; // 7 + j*5 
		#20; wea = 1; dina = 32'h000c_000a; // 12 + j*10 
		#20; wea = 1; dina = 32'h000b_0009; // 11 + j*9 
		#20; wea = 0; dina = 32'hxxxx_xxxx;
		
		// Load the instructions (only affects the raddr1, raddr0, and waddr)
		#20; inst_v = 1; rden = 0; inst = 32'h60_01_00_10; // CMPLX_MULT 
		#20; inst_v = 1; rden = 1; inst = 32'h60_03_02_11; // CMPLX_MULT 
		#20; inst_v = 1; rden = 1; inst = 32'h60_05_04_12; // CMPLX_MULT 
		#20; inst_v = 0; rden = 1; inst = 32'hxx_xx_xx_xx;
		#20; rden = 0; 
		
		// write back the 3 results generated by the ALU
        #20; wben = 1; 
        #20; wben = 1; dina = 32'h000a_000a; 
        #20; wben = 1; dina = 32'h001a_0052; 
        #20; wben = 0; dina = 32'h002a_00da; 
        #20; wben = 0; dina = 32'hxxxx_xxxx;
//        #20; inst_v = 1; rden = 0; inst = 32'h60_90_8F_13; // CMPLX_MULT 
//        #20; inst_v = 1; rden = 1; inst = 32'h60_92_91_14; // CMPLX_MULT 
//        #20; inst_v = 0; rden = 1; inst = 0;
//        #20; rden = 0;
		
		#20; web = 1; dinb = 32'h1100_1100; 
		#20; web = 1; dinb = 32'h2200_2200; 
		#20; web = 1; dinb = 32'h3300_3300; 
		#20; web = 1; dinb = 32'h4400_4400;
		#20; web = 0; dinb = 32'hxxxx_xxxx;
		#20; inst_v = 1; rden = 0; inst = 32'hxx_90_8F_xx; 
		#20; inst_v = 1; rden = 1; inst = 32'hxx_92_91_xx; 
		#20; inst_v = 0; rden = 1; inst = 32'hxx_xx_xx_xx;
		#20; rden = 0;
		
		#1000;
		
    end

endmodule
