// Data & Instructions
`define DATA_WIDTH     16
`define INST_WIDTH     64

// DSP48E2
`define PORTA_WIDTH    30
`define PORTB_WIDTH    18
`define PORTC_WIDTH    48
`define PORTP_WIDTH    48
`define ALUMODE_WIDTH   4
`define INMODE_WIDTH    5
`define OPMODE_WIDTH    7   

// Memories
`define DM_ADDR_WIDTH   8
`define IM_ADDR_WIDTH   8

// Top PE
`define PE_NUM          8
`define REG_NUM        32
`define REG_ADDR_WIDTH  5