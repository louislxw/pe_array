`define DATA_WIDTH     16
`define REG_ADDR_WIDTH  8
`define DM_ADDR_WIDTH 	8
`define IM_ADDR_WIDTH 	8
`define PORTAWIDTH     30
`define PORTBWIDTH     18
`define PORTCWIDTH     48
`define PORTPWIDTH     48